// import l1d_verif_package::*;
class l1d_downstream_trig_pkg;
    rand bit [VERIF_ADDR_WIDTH-1:0] req_addr    ;
    event                           req_trig    ;
endclass