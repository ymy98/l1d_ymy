class l1d_cfg;
    bit debug_en = 1;
endclass:l1d_cfg