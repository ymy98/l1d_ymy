module l1d_data_wr_adapter(
    input  logic clk             ,
    input  logic rst_n           ,
    input  logic downstream_rdy  ,
    output logic downstream_vld  ,
    output logic downstream_pld  
);

endmodule